module sbc_system (

);

endmodule
